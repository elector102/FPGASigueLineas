----TB
--LIBRARY ieee ;
--USE ieee.std_logic_1164.all ;
--
--Entity Tb is
--End Tb;
--
--ARCHITECTURE Behavior OF Tb IS
--
--Signal	CLK_50M :  std_logic;
--Signal	Sel_freq : std_logic_vector (2 downto 0):="000";
--Signal	Sel_cont : std_logic_vector (1 downto 0):="11";
--Signal	Up_down_0 : std_logic:='1'; -- Contador 1
--Signal	Up_down_1 : std_logic:='0'; -- Contador 2
--Signal	Areset : std_logic:='1';
--Signal	Rst_cont : std_logic:='0';
--Signal	Pll_locked : std_logic:='0';
--Signal	Out_7 : std_logic_vector (6 downto 0) :="1111111";
--
--COMPONENT pwm is
--
--generic (num_de_cont:integer := 4);
--PORT(
--        clk    : IN  STD_LOGIC;
--        reset  : IN  STD_LOGIC;
--        entrada: IN  STD_LOGIC_VECTOR(6 downto 0);
--        salida : OUT STD_LOGIC);
--END COMPONENT;
--
--BEGIN
--U1: TOP
--PORT MAP(CLK_50M, Sel_freq, Sel_cont, Up_down_0, Up_down_1, Areset, Rst_cont, Pll_locked, Out_7);
--
--Process
--	BEGIN
--	CLK_50M<='1';
--	wait for 10 ns;
--	CLK_50M<='0';
--	wait for 10 ns;
--End process;
--
--Process
--	BEGIN
--	wait until (rising_edge(Pll_locked));
--	Rst_cont <= '1';
--	Sel_freq <= "000";
--	Sel_cont <= "00";
--	wait for 1 ms;
--	Up_down_0 <='0';
--	wait for 0.6 ms;
--	Rst_cont <= '0';
--	wait for 0.2 ms;
--	Rst_cont <= '1';
--	Sel_freq <= "001";
--	Sel_cont <= "10";
--	wait for 2 ms;
--	Sel_freq <= "000";
--	Sel_cont <= "11";
--	wait for 1.2 ms; --5ms
--End process;
--
--END Behavior ;